module sign_ext
#(parameter Type_U = 7'b011_0111,
  parameter Type_J = 7'b110_1111,
  parameter Type_B = 7'b110_0011,
  parameter Type_Ijalr = 7'b110_0111,
  parameter Type_I_l = 7'b000_0011,
  parameter Type_S = 7'b010_0011,
  parameter Type_I = 7'b001_0011
)
(
	input [31:0] iv_Data,
	output [31:0] ov_Data

);

reg [31:0] ov_Data_Q;

assign ov_Data = ov_Data_Q;

always@*
begin
	case(iv_Data[6:0])
// ------------------------------ Tipo I -------------------------------------------------------------
		Type_Ijalr,Type_I_l, Type_I:
			begin
				if(iv_Data[31] == 1)
				begin
					ov_Data_Q = {20'b1111_1111_1111_1111_1111,iv_Data[31:20]};
				end
				else
				begin
					ov_Data_Q = {20'b0000_0000_0000_0000_0000,iv_Data[31:20]};
				end
			end
// ------------------------------ Tipo I -------------------------------------------------------------

// ------------------------------ Tipo S -------------------------------------------------------------		
		Type_S:
			begin
				if(iv_Data[31] == 1)
				begin
					ov_Data_Q = {20'b1111_1111_1111_1111_1111,iv_Data[31:25],iv_Data[11:7]};
				end
				else
				begin
					ov_Data_Q = {20'b0000_0000_0000_0000_0000,iv_Data[31:25],iv_Data[11:7]};
				end
			end
// ------------------------------ Tipo S -------------------------------------------------------------	

// ------------------------------ Tipo B -------------------------------------------------------------	
		Type_B: 
			begin
				if(iv_Data[31] == 1)
				begin
					ov_Data_Q = {19'b111_1111_1111_1111_1111,iv_Data[31],iv_Data[7],iv_Data[30:25],iv_Data[11:8],1'b0};
				end
				else
				begin
					ov_Data_Q = {19'b000_0000_0000_0000_0000,iv_Data[31],iv_Data[7],iv_Data[30:25],iv_Data[11:8],1'b0};
				end
			end
// ------------------------------ Tipo B -------------------------------------------------------------

// ------------------------------ Tipo U -------------------------------------------------------------	
		Type_U,7'b001_0111: ov_Data_Q = {iv_Data[31:12],12'b0};
// ------------------------------ Tipo U -------------------------------------------------------------

// ------------------------------ Tipo J -------------------------------------------------------------		
		Type_J:
			begin
				if(iv_Data[31] == 1)
				begin
					ov_Data_Q = {11'b111_1111_1111,iv_Data[31],iv_Data[19:12],iv_Data[20],iv_Data[30:21],1'b0};
				end
				else
				begin
					ov_Data_Q = {11'b000_0000_0000,iv_Data[31],iv_Data[19:12],iv_Data[20],iv_Data[30:21],1'b0};
				end
			end
// ------------------------------ Tipo J -------------------------------------------------------------
		default: ov_Data_Q = 32'b0;
	endcase
end

endmodule 