module ADD_4_Bench();

	reg i_Clk;
	reg i_Rst;
	reg i_Enb;
	reg [31:0] iv_Dir;
	wire [31:0] ov_Dir;
	
	
ADD_4 ADD_4(
	.i_Clk(i_Clk),
	.i_Rst(i_Rst),
	.i_Enb(i_Enb),
	.iv_Dir(iv_Dir),
	.ov_Dir(ov_Dir)
);


initial
begin
	i_Clk = 0;
	i_Rst = 1;
	i_Enb = 1;
	iv_Dir = 0;
	#100;
	i_Rst = 0;
	repeat(10)
	begin
		iv_Dir <= ov_Dir;
		#50;
	end
end


always
begin
	i_Clk = ~i_Clk;
	#20;
end


endmodule 